// ALU Operations
`define ALU_NOP 5'd0
`define ADD 5'd1
`define SUB 5'd2
`define XOR 5'd3
`define OR 5'd4
`define AND 5'd5
`define SLL 5'd6
`define SRL 5'd7
`define SRA 5'd8
`define SLT 5'd9
`define SLTU 5'd10
`define ADDI 5'd16
`define XORI 5'd17
`define ORI 5'd18
`define ANDI 5'd19
`define SLLI 5'd20
`define SRLI 5'd21
`define SRAI 5'd22
`define SLTI 5'd23
`define SLTIU 5'd24
`define LUI 5'd28
`define AUIPC 5'd29
