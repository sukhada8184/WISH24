module ripple_carry_adder#(
    parameter   DATA_WD=4
)(
    input   logic   [DATA_WD-1:0]   i_a,
    input   logic   [DATA_WD-1:0]   i_b,
    input   logic                   i_c,
    output  logic   [DATA_WD:0]     o_arith_out
);


    assign o_arith_out = 'b0;


endmodule
    
